module logic_design()
{

}